*** SPICE deck for cell inv_VTC{sch} from library CMOScells
*** Created on Mon Jan 15, 2024 12:06:52
*** Last revised on Mon Oct 14, 2024 23:44:25
*** Written on Thu Dec 26, 2024 12:42:01 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT CMOScells__inv FROM CELL inv{sch}
.SUBCKT CMOScells__inv a y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 y a gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd a y vdd PMOS L=0.6U W=3.6U
.ENDS CMOScells__inv

.global gnd vdd

*** TOP LEVEL CELL: inv_VTC{sch}
Xinv@0 A Y1 CMOScells__inv
Xinv@1 Y1 Y2 CMOScells__inv
Xinv@2 Y2 Y3 CMOScells__inv
Xinv@3 Y3 Y4 CMOScells__inv
Xinv@4 Y4 Y5 CMOScells__inv
Xinv@5 Y5 Y6 CMOScells__inv

* Spice Code nodes in cell cell 'inv_VTC{sch}'
.include C:\ElectricBinary\CMOScells\CMOScells\C5_models.txt
Vdd vdd 0 DC 5
Vgnd gnd 0 DC 0
Va A gnd pulse 0 5 0 0.01n 0.01n 250u 500u
.trans 0 1.5m
.END
